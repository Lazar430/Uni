module test(input [3:0]c, output f);
   f = ;
endmodule
