module hex(input [3 : 0]c, output [6:0]seg);
   assign seg[6] = ( ~(c[3]) & ~(c[2]) & ~(c[1]) & (c[0]) ) |
	    ( (c[3]) & ~(c[2]) & ~(c[1]) & ~(c[0]) ) |
	    ( (c[3]) & (c[2]) & ~(c[1]) & (c[0]) ) |
	    ( (c[3]) & ~(c[2]) & (c[1]) & (c[0]) );

   assign seg[5] = ( (c[3]) & (c[1]) & (c[0]) ) |
	    ( (c[3]) & (c[2]) & ~(c[0]) ) |
	    ( (c[2]) & (c[1]) & ~(c[0]) );

   assign seg[4] = ( ~(c[3]) & ~(c[2]) & ~(c[1]) & ~(c[0]) ) |
	    ( (c[3]) & (c[2]) & (c[1])) |
	    ( (c[3]) & (c[2]) & ~(c[0]) );

   assign seg[3] = ( (c[2]) & (c[1]) & (c[0]) ) |
	    ( ~(c[3]) & ~(c[2]) & ~(c[1]) & (c[0]) ) |
	    ( ~(c[3]) & (c[2]) & ~(c[1]) & (c[0]) ) |
	    ( ~(c[3]) & (c[2]) & ~(c[1]) & ~(c[0]) );

   assign seg[2] = ( ~(c[3]) & (c[2]) & ~(c[1]) ) |
	    ( ~(c[3]) & (c[1]) & (c[0]) ) |
	    ( (c[2]) & ~(c[1]) & (c[0]) );

   assign seg[1] = ( ~(c[3]) & ~(c[2]) & (c[0]) ) |
	    ( (c[3]) & ~(c[2]) & (c[1]) ) |
	    ( (c[3]) & (c[2]) & ~(c[1]) & (c[0]) );

   assign seg[0] = ( ~(c[3]) & (c[2]) & (c[1]) & (c[0]) ) |
	    ( ~(c[3]) & ~(c[2]) & ~(c[1]) ) |
	    ( (c[3]) & (c[2]) & ~(c[1]) & ~(c[0]) );
   
endmodule // hex
