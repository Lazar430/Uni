module hex(input [3 : 0]i, output [6:0]seg);
   assign seg[6] = ( ~(i[3]) & (i[2]) & ~(i[1]) & (i[0]) ) |
		   ( ~(i[3]) & ~(i[2]) & (i[1]) & (i[0]) ) |
		   ( ~(i[3]) & (i[2]) & (i[1]) & (i[0]) ) |
		   ( (i[3]) & (i[2]) & (i[1]) & ~(i[0]) );

   assign seg[5] = ( ~(i[3]) & (i[2]) & ~(i[1]) & (i[0]) ) |
		   ( ~(i[2]) & (i[1]) & (i[0]) ) |
		   ( (i[3]) & (i[2]) & (i[1]) ) |
		   ( (i[3]) & ~(i[2]) & (i[0]) );

   assign seg[4] = ( (i[3]) & ~(i[2]) & ~(i[1]) & ~(i[0]) ) |
		   ( (i[3]) & (i[1]) & (i[0]) ) |
		   ( ~(i[2]) & (i[1]) & (i[0]) );
   

   assign seg[3] = ( ~(i[3]) & (i[2]) & ~(i[1]) & ~(i[0]) ) |
		   ( ~(i[3]) & ~(i[2]) & ~(i[1]) & (i[0]) ) |
		   ( (i[3]) & (i[2]) & (i[1]) ) |
		   ( (i[3]) & ~(i[2]) & (i[1]) & ~(i[0]) );

   assign seg[2] = ( (i[2]) & ~(i[1]) ) |
		   ( ~(i[3]) & ~(i[1]) & (i[0]) ) |
		   ( ~(i[3]) & (i[2]) & ~(i[1]) );

   assign seg[1] = ( ~(i[3]) & (i[2]) & (i[1]) & (i[0]) ) |
		   ( (i[2]) & ~(i[1]) & ~(i[0]) ) |
		   ( (i[3]) & ~(i[1]) & ~(i[0]) ) |
		   ( (i[3]) & (i[2]) & (i[1]) );

   assign seg[0] = ( (i[3]) & (i[2]) & ~(i[1]) & (i[0]) ) |
		   ( ~(i[3]) & ~(i[1]) & ~(i[0]) );
   
endmodule // hex
